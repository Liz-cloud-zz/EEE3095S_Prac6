// Code your testbench here
// or browse Examples
`include "tb_simple_CPU.v"